// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

// Wrapper for a cv32e40p core and optional FPU
// Contributor: Davide Schiavone <davide@openhwgroup.org>

module cv32e40p_wrapper
#(
    parameter PULP_XPULP       = 0, // PULP ISA Extension (incl. custom CSRs and hardware loop, excl. p.elw)
    parameter PULP_CLUSTER     = 0, // PULP Cluster interface (incl. p.elw)
    parameter FPU              = 0, // Floating Point Unit (interfaced via APU interface)
    parameter PULP_ZFINX       = 0, // Float-in-General Purpose registers
    parameter NUM_MHPMCOUNTERS = 1
) (
    // Clock and Reset
    input logic clk_i,
    input logic rst_ni,

    input logic pulp_clock_en_i,  // PULP clock enable (only used if PULP_CLUSTER = 1)
    input logic scan_cg_en_i,  // Enable all clock gates for testing

    // Core ID, Cluster ID, debug mode halt address and boot address are considered more or less static
    input logic [31:0] boot_addr_i,
    input logic [31:0] mtvec_addr_i,
    input logic [31:0] dm_halt_addr_i,
    input logic [31:0] hart_id_i,
    input logic [31:0] dm_exception_addr_i,

    // Instruction memory interface
    output logic        instr_req_o,
    input  logic        instr_gnt_i,
    input  logic        instr_rvalid_i,
    output logic [31:0] instr_addr_o,
    input  logic [31:0] instr_rdata_i,

    // Data memory interface
    output logic        data_req_o,
    input  logic        data_gnt_i,
    input  logic        data_rvalid_i,
    output logic        data_we_o,
    output logic [ 3:0] data_be_o,
    output logic [31:0] data_addr_o,
    output logic [31:0] data_wdata_o,
    input  logic [31:0] data_rdata_i,

    // Interrupt inputs
    input  logic [31:0] irq_i,  // CLINT interrupts + CLINT extension interrupts
    output logic        irq_ack_o,
    output logic [ 4:0] irq_id_o,

    // Debug Interface
    input  logic debug_req_i,
    output logic debug_havereset_o,
    output logic debug_running_o,
    output logic debug_halted_o,

    // CPU Control Signals
    input  logic fetch_enable_i,
    output logic core_sleep_o
);
 
  import cv32e40p_apu_core_pkg::*;

  // Core to FPU
  logic                               apu_req;
  logic [    APU_NARGS_CPU-1:0][31:0] apu_operands;
  logic [      APU_WOP_CPU-1:0]       apu_op;
  logic [ APU_NDSFLAGS_CPU-1:0]       apu_flags;

  // FPU to Core
  logic                               apu_gnt;
  logic                               apu_rvalid;
  logic [                 31:0]       apu_rdata;
  logic [ APU_NUSFLAGS_CPU-1:0]       apu_rflags;

  // Instantiate the Core
  cv32e40p_core #(
    .PULP_XPULP      (PULP_XPULP),
    .PULP_CLUSTER    (PULP_CLUSTER),
    .FPU             (FPU),
    .PULP_ZFINX      (PULP_ZFINX),
    .NUM_MHPMCOUNTERS(NUM_MHPMCOUNTERS)
  ) core_i (
    .clk_i               (clk_i              ),
    .rst_ni              (rst_ni             ),

    .pulp_clock_en_i     (pulp_clock_en_i    ),
    .scan_cg_en_i        (scan_cg_en_i       ),

    .boot_addr_i         (boot_addr_i        ),
    .mtvec_addr_i        (mtvec_addr_i       ),
    .dm_halt_addr_i      (dm_halt_addr_i     ),
    .hart_id_i           (hart_id_i          ),
    .dm_exception_addr_i (dm_exception_addr_i),

    .instr_req_o         (instr_req_o        ),
    .instr_gnt_i         (instr_gnt_i        ),
    .instr_rvalid_i      (instr_rvalid_i     ),
    .instr_addr_o        (instr_addr_o       ),
    .instr_rdata_i       (instr_rdata_i      ),

    .data_req_o          (data_req_o         ),
    .data_gnt_i          (data_gnt_i         ),
    .data_rvalid_i       (data_rvalid_i      ),
    .data_we_o           (data_we_o          ),
    .data_be_o           (data_be_o          ),
    .data_addr_o         (data_addr_o        ),
    .data_wdata_o        (data_wdata_o       ),
    .data_rdata_i        (data_rdata_i       ),

    .apu_req_o           (apu_req            ),
    .apu_gnt_i           (apu_gnt            ),
    .apu_operands_o      (apu_operands       ),
    .apu_op_o            (apu_op             ),
    .apu_flags_o         (apu_flags          ),
    .apu_rvalid_i        (apu_rvalid         ),
    .apu_result_i        (apu_rdata          ),
    .apu_flags_i         (apu_rflags         ),

    .irq_i               (irq_i              ),
    .irq_ack_o           (irq_ack_o          ),
    .irq_id_o            (irq_id_o           ),

    .debug_req_i         (debug_req_i        ),
    .debug_havereset_o   (debug_havereset_o  ),
    .debug_running_o     (debug_running_o    ),
    .debug_halted_o      (debug_halted_o     ),

    .fetch_enable_i      (fetch_enable_i     ),
    .core_sleep_o        (core_sleep_o       )
  );

  generate
    if (FPU) begin : fpu_gen
      // Instantiate the FPU wrapper
      cv32e40p_fp_wrapper fp_wrapper_i (
        .clk_i          ( clk_i        ),
        .rst_ni         ( rst_ni       ),
        .apu_req_i      ( apu_req      ),
        .apu_gnt_o      ( apu_gnt      ),
        .apu_operands_i ( apu_operands ),
        .apu_op_i       ( apu_op       ),
        .apu_flags_i    ( apu_flags    ),
        .apu_rvalid_o   ( apu_rvalid   ),
        .apu_rdata_o    ( apu_rdata    ),
        .apu_rflags_o   ( apu_rflags    )
      );
    end else begin : no_fpu_gen
      // Drive FPU output signals to 0
      assign apu_gnt    = '0;
      assign apu_rvalid = '0;
      assign apu_rdata  = '0;
      assign apu_rflags = '0;
    end
  endgenerate

endmodule
