// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

/////////////////////////////////////////////////////////////////////////////////////////////////
//                                                                                             //
// Author:                        Francesco Minervini - minervif@student.ethz.ch               //
//                                                                                             //
// Additional contributions by:                                                                //
//                                                                                             //
// Design Name:                   Top level module including riscv core and perturbation       //
//                                module                                                       //
// Project Name:                  TB RISC-V                                                    //
// Language:                      SystemVerilog                                                //
//                                                                                             //
// Description:                   This module is instantiated in the core_region.sv code       //
//                                when the parameter TB_RISCV is set to 1.                     //
//                                This module instantiates one between zero_riscy or riscy     //
//                                core depending on the value of USE_ZERO_RISCY, then          //
//                                it also instantiates and connects the core to the            //
//                                perturbation module.                                         //
//                                                                                             //
/////////////////////////////////////////////////////////////////////////////////////////////////

module tb_cv32e40p_core
#(
  parameter INSTR_RDATA_WIDTH   = 32,
  parameter WAPUTYPE            =  0,
  parameter APU_NARGS_CPU       =  3,
  parameter APU_WOP_CPU         =  6,
  parameter APU_NDSFLAGS_CPU    = 15,
  parameter APU_NUSFLAGS_CPU    =  5,
  parameter SIMCHECKER          =  0,
  parameter PULP_CLUSTER        =  0,
  parameter FPU                 =  0,
  parameter PULP_ZFINX          =  0,
  parameter DM_HALTADDRESS      = 32'h1A110800
)
(
  // Clock and Reset
  input  logic        clk_i,
  input  logic        rst_ni,

  input  logic        clock_en_i,    // enable clock, otherwise it is gated
  input  logic        test_en_i,     // enable all clock gates for testing

  input  logic        fregfile_disable_i,  // disable the fp regfile, using int regfile instead

  // Core ID, Cluster ID and boot address are considered more or less static
  input  logic [31:0] boot_addr_i,
  input  logic [ 3:0] core_id_i,
  input  logic [ 5:0] cluster_id_i,

  // Instruction memory interface
  output logic                         instr_req_o,
  input  logic                         instr_gnt_i,
  input  logic                         instr_rvalid_i,
  output logic                  [31:0] instr_addr_o,
  input  logic [INSTR_RDATA_WIDTH-1:0] instr_rdata_i,

  // Data memory interface
  output logic        data_req_o,
  input  logic        data_gnt_i,
  input  logic        data_rvalid_i,
  output logic        data_we_o,
  output logic [3:0]  data_be_o,
  output logic [31:0] data_addr_o,
  output logic [31:0] data_wdata_o,
  input  logic [31:0] data_rdata_i,
  // apu-interconnect
  // handshake signals
  output logic                       apu_master_req_o,
  output logic                       apu_master_ready_o,
  input logic                        apu_master_gnt_i,
  // request channel
  output logic [31:0]                 apu_master_operands_o [APU_NARGS_CPU-1:0],
  output logic [APU_WOP_CPU-1:0]      apu_master_op_o,
  output logic [WAPUTYPE-1:0]         apu_master_type_o,
  output logic [APU_NDSFLAGS_CPU-1:0] apu_master_flags_o,
  // response channel
  input logic                        apu_master_valid_i,
  input logic [31:0]                 apu_master_result_i,
  input logic [APU_NUSFLAGS_CPU-1:0] apu_master_flags_i,

  // Interrupt inputs
  input  logic        irq_i,                 // level sensitive IR lines
  input  logic [4:0]  irq_id_i,
  output logic        irq_ack_o,
  output logic [4:0]  irq_id_o,

  // Debug Interface
  input  logic        debug_req_i,
  output logic        debug_gnt_o,
  output logic        debug_rvalid_o,
  input  logic [14:0] debug_addr_i,
  input  logic        debug_we_i,
  input  logic [31:0] debug_wdata_i,
  output logic [31:0] debug_rdata_o,
  output logic        debug_halted_o,
  input  logic        debug_halt_i,
  input  logic        debug_resume_i,

  // CPU Control Signals
  input  logic        fetch_enable_i,
  output logic        core_busy_o
);

localparam PERT_REGS = 15;

//////////////////////////////////////////////////////////////
//Internal signals to connect core and perturbation module
/////////////////////////////////////////////////////////////

// Additional instruction signals

logic                          instr_req_int;
logic                          instr_grant_int;
logic                          instr_rvalid_int;
logic [31:0]                   instr_addr_int;
logic [INSTR_RDATA_WIDTH-1:0]  instr_rdata_int;

// Additional data signals
logic                          data_req_int;
logic                          data_grant_int;
logic                          data_rvalid_int;
logic                          data_we_int;
logic [3:0]                    data_be_int;
logic [31:0]                   data_addr_int;
logic [31:0]                   data_wdata_int;
logic [31:0]                   data_rdata_int;

// Additional signals for pertubation/debug registers
logic                          debug_req_int;
logic                          debug_grant_int;
logic                          debug_rvalid_int;
logic                          debug_we_int;
logic [14:0]                   debug_addr_int;
logic [31:0]                   debug_wdata_int;
logic [31:0]                   debug_rdata_int;

// Additional interrupt signals
logic                          irq_int;
logic                          irq_ack_int;
logic [4:0]                    irq_id_int;
logic [4:0]                    irq_core_resp_id_int;



  cv32e40p_core
  #(
    .PULP_CLUSTER(PULP_CLUSTER),
    .FPU(FPU),
    .PULP_ZFINX(PULP_ZFINX),
    .DM_HALTADDRESS(DM_HALTADDRESS)
    )
  core_i
  (
    .clk_i                          ( clk_i                   ),
    .rst_ni                         ( rst_ni                  ),

    .clock_en_i                     ( clock_en_i              ),
    .test_en_i                      ( test_en_i               ),

    .boot_addr_i                    ( boot_addr_i             ),
    .core_id_i                      ( core_id_i               ),
    .cluster_id_i                   ( cluster_id_i            ),

    .instr_req_o                    ( instr_req_int           ),
    .instr_gnt_i                    ( instr_grant_int         ),
    .instr_rvalid_i                 ( instr_rvalid_int        ),
    .instr_addr_o                   ( instr_addr_int          ),
    .instr_rdata_i                  ( instr_rdata_int         ),

    .data_req_o                     ( data_req_int            ),
    .data_gnt_i                     ( data_grant_int          ),
    .data_rvalid_i                  ( data_rvalid_int         ),
    .data_we_o                      ( data_we_int             ),
    .data_be_o                      ( data_be_int             ),
    .data_addr_o                    ( data_addr_int           ),
    .data_wdata_o                   ( data_wdata_int          ),
    .data_rdata_i                   ( data_rdata_int          ),

    .apu_master_req_o               ( apu_master_req_o        ),
    .apu_master_ready_o             ( apu_master_ready_o      ),
    .apu_master_gnt_i               ( apu_master_gnt_i        ),
    .apu_master_operands_o          ( apu_master_operands_o   ),
    .apu_master_op_o                ( apu_master_op_o         ),
    .apu_master_type_o              ( apu_master_type_o       ),
    .apu_master_flags_o             ( apu_master_flags_o      ),
    .apu_master_valid_i             ( apu_master_valid_i      ),
    .apu_master_result_i            ( apu_master_result_i     ),
    .apu_master_flags_i             ( apu_master_flags_i      ),

    .irq_software_i                 ( 1'b0                    ),
    .irq_timer_i                    ( 1'b0                    ), 
    .irq_external_i                 ( 1'b0                    ), 
    .irq_fast_i                     ( 15'b0                   ), 
    .irq_nmi_i                      ( 1'b0                    ), 
    .irq_fastx_i                    ( 32'b0                   ), 
    .irq_ack_o                      ( irq_ack_int             ), 
    .irq_id_o                       ( irq_core_resp_id_int    ), 

    .debug_req_i                    ( debug_req_int           ),

    .fetch_enable_i                 ( fetch_enable_i          ),
    .core_busy_o                    ( core_busy_o             ),

    .fregfile_disable_i             ( fregfile_disable_i      )
  );

  // Perturbation module instance
  cv32e40p_perturbation
  #(
   .PERT_REGS                      ( PERT_REGS         ),
   .INSTR_RDATA_WIDTH              ( INSTR_RDATA_WIDTH )
  )
  perturbation_i
  (
    .clk_i                         ( clk_i                  ),
    .rst_ni                        ( rst_ni                 ),

    .pert_instr_req_i              ( instr_req_int          ),
    .pert_instr_req_o              ( instr_req_o            ),
    .pert_instr_grant_i            ( instr_gnt_i            ),
    .pert_instr_grant_o            ( instr_grant_int        ),
    .pert_instr_rvalid_i           ( instr_rvalid_i         ),
    .pert_instr_rvalid_o           ( instr_rvalid_int       ),
    .pert_instr_addr_i             ( instr_addr_int         ),
    .pert_instr_addr_o             ( instr_addr_o           ),
    .pert_instr_rdata_i            ( instr_rdata_i          ),
    .pert_instr_rdata_o            ( instr_rdata_int        ),

    .pert_data_req_i               ( data_req_int           ),
    .pert_data_req_o               ( data_req_o             ),
    .pert_data_grant_i             ( data_gnt_i             ),
    .pert_data_grant_o             ( data_grant_int         ),
    .pert_data_rvalid_i            ( data_rvalid_i          ),
    .pert_data_rvalid_o            ( data_rvalid_int        ),
    .pert_data_we_i                ( data_we_int            ),
    .pert_data_we_o                ( data_we_o              ),
    .pert_data_be_i                ( data_be_int            ),
    .pert_data_be_o                ( data_be_o              ),
    .pert_data_addr_i              ( data_addr_int          ),
    .pert_data_addr_o              ( data_addr_o            ),
    .pert_data_wdata_i             ( data_wdata_int         ),
    .pert_data_wdata_o             ( data_wdata_o           ),
    .pert_data_rdata_i             ( data_rdata_i           ),
    .pert_data_rdata_o             ( data_rdata_int         ),

    .pert_debug_req_i              ( debug_req_i            ),
    .pert_debug_req_o              ( debug_req_int          ),
    .pert_debug_gnt_i              ( debug_grant_int        ),
    .pert_debug_gnt_o              ( debug_gnt_o            ),
    .pert_debug_rvalid_i           ( debug_rvalid_int       ),
    .pert_debug_rvalid_o           ( debug_rvalid_o         ),
    .pert_debug_we_i               ( debug_we_i             ),
    .pert_debug_we_o               ( debug_we_int           ),
    .pert_debug_addr_i             ( debug_addr_i           ),
    .pert_debug_addr_o             ( debug_addr_int         ),
    .pert_debug_wdata_i            ( debug_wdata_i          ),
    .pert_debug_wdata_o            ( debug_wdata_int        ),
    .pert_debug_rdata_i            ( debug_rdata_int        ),
    .pert_debug_rdata_o            ( debug_rdata_o          ),

    .pert_irq_i                    ( irq_i                  ),
    .pert_irq_o                    ( irq_int                ),
    .pert_irq_id_i                 ( irq_id_i               ),
    .pert_irq_id_o                 ( irq_id_int             ),
    .pert_irq_ack_i                ( irq_ack_int            ),
    .pert_irq_ack_o                ( irq_ack_o              ),
    .pert_irq_core_resp_id_i       ( irq_core_resp_id_int   ),
    .pert_irq_core_resp_id_o       ( irq_id_o               ),
    .pert_pc_id_i                  ( core_i.pc_id           )
  );


   `ifndef VERILATOR
   generate
       if(SIMCHECKER) begin: ri5cy_simchecker
          cv32e40p_simchecker simchecker_i
          (
            .clk              ( core_i.clk_i                                ),
            .rst_n            ( core_i.rst_ni                               ),

            .fetch_enable     ( core_i.fetch_enable_i                       ),
            .boot_addr        ( core_i.boot_addr_i                          ),
            .core_id          ( core_i.core_id_i                            ),
            .cluster_id       ( core_i.cluster_id_i                         ),

            .instr_compressed ( core_i.if_stage_i.fetch_rdata[15:0]         ),
            .if_valid         ( core_i.if_stage_i.if_valid                  ),
            .pc_set           ( core_i.pc_set                               ),


            .pc               ( core_i.id_stage_i.pc_id_i                   ),
            .instr            ( core_i.id_stage_i.instr                     ),
            .is_compressed    ( core_i.is_compressed_id                     ),
            .id_valid         ( core_i.id_stage_i.id_valid_o                ),
            .is_decoding      ( core_i.id_stage_i.is_decoding_o             ),
            .is_illegal       ( core_i.id_stage_i.illegal_insn_dec          ),
            .is_interrupt     ( core_i.is_interrupt                         ),
            .irq_no           ( core_i.irq_id_i                             ),
            .pipe_flush       ( core_i.id_stage_i.controller_i.pipe_flush_i ),
            .irq_i            ( core_i.irq_i                                ),
            .is_mret          ( core_i.id_stage_i.controller_i.mret_insn_i  ),

            .int_enable       ( core_i.id_stage_i.m_irq_enable_i            ),

            .lsu_ready_wb     ( core_i.lsu_ready_wb                         ),
            .apu_ready_wb     ( core_i.apu_ready_wb                         ),
            .wb_contention    ( core_i.ex_stage_i.wb_contention             ),

            .apu_en_id        ( core_i.id_stage_i.apu_en                    ),
            .apu_req          ( core_i.ex_stage_i.apu_req                   ),
            .apu_gnt          ( core_i.ex_stage_i.apu_gnt                   ),
            .apu_valid        ( core_i.ex_stage_i.apu_valid                 ),
            .apu_singlecycle  ( core_i.ex_stage_i.apu_singlecycle           ),
            .apu_multicycle   ( core_i.ex_stage_i.apu_multicycle            ),
            .apu_latency      ( core_i.ex_stage_i.apu_lat_i                 ),
            .apu_active       ( core_i.ex_stage_i.apu_active                ),
            .apu_en_ex        ( core_i.ex_stage_i.apu_en_i                  ),

            .ex_valid         ( core_i.ex_valid                             ),
            .ex_reg_addr      ( core_i.id_stage_i.registers_i.waddr_b_i     ),

            .ex_reg_we        ( core_i.id_stage_i.registers_i.we_b_i        ),
            .ex_reg_wdata     ( core_i.id_stage_i.registers_i.wdata_b_i     ),

            .ex_data_req      ( core_i.data_req_o                           ),
            .ex_data_gnt      ( core_i.data_gnt_i                           ),
            .ex_data_we       ( core_i.data_we_o                            ),
            .ex_data_addr     ( core_i.data_addr_o                          ),
            .ex_data_wdata    ( core_i.data_wdata_o                         ),

            .lsu_misaligned   ( core_i.data_misaligned                      ),
            .wb_bypass        ( core_i.ex_stage_i.branch_in_ex_i            ),

            .wb_valid         ( core_i.wb_valid                             ),
            .wb_reg_addr      ( core_i.id_stage_i.registers_i.waddr_a_i     ),
            .wb_reg_we        ( core_i.id_stage_i.registers_i.we_a_i        ),
            .wb_reg_wdata     ( core_i.id_stage_i.registers_i.wdata_a_i     ),
            .wb_data_rvalid   ( core_i.data_rvalid_i                        ),
            .wb_data_rdata    ( core_i.data_rdata_i                         )
          );
        end
   endgenerate
   `endif

endmodule // tb_cv32e40p_core
