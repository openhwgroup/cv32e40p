///////////////////////////////////////////////////////////////////////////////
//                                                                           //
// RISC-V Checker                                                            //
//                                                                           //
// This material contains trade secrets or otherwise confidential            //
// information owned by Siemens Industry Software Inc. or its affiliates     //
// (collectively, "SISW"), or its licensors. Access to and use of this       //
// information is strictly limited as set forth in the Customer's applicable //
// agreements with SISW.                                                     //
//                                                                           //
// This material may not be copied, distributed, or otherwise disclosed      //
// outside of the Customer's facilities without the express written          //
// permission of SISW, and may not be used in any way not expressly          //
// authorized by SISW.                                                       //
//                                                                           //
///////////////////////////////////////////////////////////////////////////////




This file is available only to Siemens EDA OneSpin customers and is available by submitting a request to Siemens support center to get it.
